library ieee;
use ieee.std_logic_1164.all;

entity practica_1 is
	port (y: in std_logic_vector(3 downto 0);
 	z: out std_logic_vector(3 downto 0));
end practica_1;
